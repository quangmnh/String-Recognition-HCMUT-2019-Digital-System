module quads1(qout,qin);
	output reg qout;
	input qin;
endmodule 